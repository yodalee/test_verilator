package pkg;

typedef logic [4:0] qbit;

endpackage