`include "pkg.sv"

module sub ();
endmodule