`include "sub.sv"
`include "pkg.sv"

import pkg::*;

module top ();

sub i_sub();

endmodule